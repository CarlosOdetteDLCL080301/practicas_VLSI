library ieee;
use ieee.std_logic_1164.all;

entity ControlTREN is
	port(
	
	);
end entity;

architecture arq_ControlTREN of ControlTREN is

end architecture;